library verilog;
use verilog.vl_types.all;
entity L1P3_vlg_vec_tst is
end L1P3_vlg_vec_tst;
