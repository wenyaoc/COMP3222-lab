library verilog;
use verilog.vl_types.all;
entity L9P1board_vlg_vec_tst is
end L9P1board_vlg_vec_tst;
