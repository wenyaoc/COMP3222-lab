library verilog;
use verilog.vl_types.all;
entity L3P4_vlg_vec_tst is
end L3P4_vlg_vec_tst;
