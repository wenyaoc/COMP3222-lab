library verilog;
use verilog.vl_types.all;
entity L9P2_vlg_vec_tst is
end L9P2_vlg_vec_tst;
