library verilog;
use verilog.vl_types.all;
entity L3P2 is
    port(
        Clk             : in     vl_logic;
        D               : in     vl_logic;
        Q               : out    vl_logic
    );
end L3P2;
