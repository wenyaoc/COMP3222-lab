library verilog;
use verilog.vl_types.all;
entity L7P2_vlg_vec_tst is
end L7P2_vlg_vec_tst;
