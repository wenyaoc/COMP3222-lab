library verilog;
use verilog.vl_types.all;
entity L1P4_vlg_vec_tst is
end L1P4_vlg_vec_tst;
