library verilog;
use verilog.vl_types.all;
entity L3P1_vlg_vec_tst is
end L3P1_vlg_vec_tst;
