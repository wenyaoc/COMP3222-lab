library verilog;
use verilog.vl_types.all;
entity L11P2_vlg_vec_tst is
end L11P2_vlg_vec_tst;
